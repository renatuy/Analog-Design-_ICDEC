magic
tech sky130A
magscale 1 2
timestamp 1729062773
<< viali >>
rect 133 1053 1140 1095
rect 133 32 1140 74
<< metal1 >>
rect 121 1095 1152 1101
rect 121 1053 133 1095
rect 1140 1053 1152 1095
rect 121 1047 1152 1053
rect 174 533 184 585
rect 236 533 246 585
rect 280 544 643 577
rect 704 542 1067 575
rect 1120 533 1130 585
rect 1182 533 1192 585
rect 121 74 1152 80
rect 121 32 133 74
rect 1140 32 1152 74
rect 121 26 1152 32
<< via1 >>
rect 184 533 236 585
rect 1130 533 1182 585
<< metal2 >>
rect 184 587 236 595
rect 1130 587 1182 595
rect 180 585 1183 587
rect 180 533 184 585
rect 236 533 1130 585
rect 1182 533 1183 585
rect 184 523 236 533
rect 1130 523 1182 533
use inverter  x1
timestamp 1728981621
transform 1 0 182 0 1 566
box -182 -566 240 562
use inverter  x2
timestamp 1728981621
transform 1 0 604 0 1 566
box -182 -566 240 562
use inverter  x3
timestamp 1728981621
transform 1 0 1026 0 1 566
box -182 -566 240 562
<< labels >>
flabel viali 361 1068 361 1068 0 FreeSans 160 0 0 0 vdd
port 3 nsew
flabel viali 365 42 365 42 0 FreeSans 160 0 0 0 gnd
port 5 nsew
flabel metal2 848 558 848 558 0 FreeSans 160 0 0 0 out
port 7 nsew
<< end >>
