magic
tech sky130A
magscale 1 2
timestamp 1729049424
<< checkpaint >>
rect -997 -2043 1945 1097
<< error_s >>
rect -51 -579 -36 -217
rect 76 -230 134 -224
rect -17 -545 -2 -251
rect 76 -264 88 -230
rect 113 -264 134 -230
rect 76 -270 134 -264
rect 10 -283 17 -273
rect 141 -283 162 -196
rect 10 -285 23 -283
rect 6 -340 23 -285
rect 141 -291 175 -283
rect 44 -311 51 -307
rect 38 -323 51 -311
rect 126 -319 172 -311
rect 38 -340 55 -323
rect 6 -537 17 -340
rect 44 -499 55 -340
rect 155 -433 172 -319
rect 183 -405 200 -340
rect 44 -515 51 -499
rect 10 -545 17 -537
rect 76 -558 134 -552
rect 76 -592 88 -558
rect 76 -598 134 -592
<< viali >>
rect -17 19 17 321
rect -17 -545 17 -251
<< metal1 >>
rect -23 321 23 333
rect -23 19 -17 321
rect 17 295 23 321
rect 17 117 132 295
rect 180 123 267 173
rect 17 19 23 117
rect -23 7 23 19
rect -23 -251 23 -239
rect -23 -545 -17 -251
rect 17 -340 23 -251
rect 141 -291 175 59
rect 217 -340 267 123
rect 17 -517 132 -340
rect 183 -405 268 -340
rect 17 -545 23 -517
rect -23 -557 23 -545
use sky130_fd_pr__pfet_01v8_XGS3BL  XM1
timestamp 0
transform 1 0 105 0 1 -411
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 0
transform 1 0 474 0 1 -473
box -211 -310 211 310
<< labels >>
flabel metal1 43 182 43 182 0 FreeSans 160 0 0 0 vdd
port 1 nsew
flabel metal1 37 -440 37 -437 0 FreeSans 160 0 0 0 gnd
port 3 nsew
flabel metal1 155 -127 155 -127 0 FreeSans 160 0 0 0 in
port 5 nsew
flabel metal1 235 -133 235 -133 0 FreeSans 160 0 0 0 out
port 7 nsew
<< end >>
